library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity FrequencyGenerator is
port(Resetn: in std_logic;
	  Clk: in std_logic;
     BPM: in std_logic_vector(10 downto 0);
	  Compas: in std_logic_vector(3 downto 0);
	  Secuencia_leds: out std_logic_vector(2 downto 0);
	  Secuencia_sonido: out std_logic);
end FrequencyGenerator;

architecture Solucion of FrequencyGenerator is
constant t_10ms: integer:= 500000;
shared variable BPM_integer: integer:= to_integer(unsigned(BPM));
shared variable freq: integer:= 0;
signal counter: std_logic_vector(26 downto 0);

begin

process(Resetn)
begin
	if Resetn='0' then freq:= 0;
	else
		case BPM_integer is
			when 30=> freq:= 100000000;
			when 31=> freq:= 96774193;
			when 32=> freq:= 93750000;
			when 33=> freq:= 90909090;
			when 34=> freq:= 88235294;
			when 35=> freq:= 85714285;
			when 36=> freq:= 83333333;
			when 37=> freq:= 81081081;
			when 38=> freq:= 78947368;
			when 39=> freq:= 76923076;
			when 40=> freq:= 75000000;
			when 41=> freq:= 73170731;
			when 42=> freq:= 71428571;
			when 43=> freq:= 69767441;
			when 44=> freq:= 68181818;
			when 45=> freq:= 66666666;
			when 46=> freq:= 65217391;
			when 47=> freq:= 63829787;
			when 48=> freq:= 62500000;
			when 49=> freq:= 61224489;
			when 50=> freq:= 60000000;
			when 51=> freq:= 58823529;
			when 52=> freq:= 57692307;
			when 53=> freq:= 56603773;
			when 54=> freq:= 55555555;
			when 55=> freq:= 54545454;
			when 56=> freq:= 53571428;
			when 57=> freq:= 52631578;
			when 58=> freq:= 51724137;
			when 59=> freq:= 50847457;
			when 60=> freq:= 50000000;
			when 61=> freq:= 49180327;
			when 62=> freq:= 48387096;
			when 63=> freq:= 47619047;
			when 64=> freq:= 46875000;
			when 65=> freq:= 46153846;
			when 66=> freq:= 45454545;
			when 67=> freq:= 44776119;
			when 68=> freq:= 44117647;
			when 69=> freq:= 43478260;
			when 70=> freq:= 42857142;
			when 71=> freq:= 42253521;
			when 72=> freq:= 41666666;
			when 73=> freq:= 41095890;
			when 74=> freq:= 40540540;
			when 75=> freq:= 40000000;
			when 76=> freq:= 39473684;
			when 77=> freq:= 38961039;
			when 78=> freq:= 38461538;
			when 79=> freq:= 37974683;
			when 80=> freq:= 37500000;
			when 81=> freq:= 37037037;
			when 82=> freq:= 36585365;
			when 83=> freq:= 36144578;
			when 84=> freq:= 35714285;
			when 85=> freq:= 35294117;
			when 86=> freq:= 34883720;
			when 87=> freq:= 34482758;
			when 88=> freq:= 34090909;
			when 89=> freq:= 33707865;
			when 90=> freq:= 33333333;
			when 91=> freq:= 32967033;
			when 92=> freq:= 32608695;
			when 93=> freq:= 32258064;
			when 94=> freq:= 31914893;
			when 95=> freq:= 31578947;
			when 96=> freq:= 31250000;
			when 97=> freq:= 30927835;
			when 98=> freq:= 30612244;
			when 99=> freq:= 30303030;
			when 100=> freq:= 30000000;
			when 101=> freq:= 29702970;
			when 102=> freq:= 29411764;
			when 103=> freq:= 29126213;
			when 104=> freq:= 28846153;
			when 105=> freq:= 28571428;
			when 106=> freq:= 28301886;
			when 107=> freq:= 28037383;
			when 108=> freq:= 27777777;
			when 109=> freq:= 27522935;
			when 110=> freq:= 27272727;
			when 111=> freq:= 27027027;
			when 112=> freq:= 26785714;
			when 113=> freq:= 26548672;
			when 114=> freq:= 26315789;
			when 115=> freq:= 26086956;
			when 116=> freq:= 25862069;
			when 117=> freq:= 25641025;
			when 118=> freq:= 25423728;
			when 119=> freq:= 25210084;
			when 120=> freq:= 25000000;
			when 121=> freq:= 24793388;
			when 122=> freq:= 24590163;
			when 123=> freq:= 24390243;
			when 124=> freq:= 24193548;
			when 125=> freq:= 24000000;
			when 126=> freq:= 23809523;
			when 127=> freq:= 23622047;
			when 128=> freq:= 23437500;
			when 129=> freq:= 23255814;
			when 130=> freq:= 23076923;
			when 131=> freq:= 22900763;
			when 132=> freq:= 22727272;
			when 133=> freq:= 22556391;
			when 134=> freq:= 22388059;
			when 135=> freq:= 22222222;
			when 136=> freq:= 22058823;
			when 137=> freq:= 21897810;
			when 138=> freq:= 21739130;
			when 139=> freq:= 21582733;
			when 140=> freq:= 21428571;
			when 141=> freq:= 21276595;
			when 142=> freq:= 21126760;
			when 143=> freq:= 20979021;
			when 144=> freq:= 20833333;
			when 145=> freq:= 20689655;
			when 146=> freq:= 20547945;
			when 147=> freq:= 20408163;
			when 148=> freq:= 20270270;
			when 149=> freq:= 20134228;
			when 150=> freq:= 20000000;
			when 151=> freq:= 19867549;
			when 152=> freq:= 19736842;
			when 153=> freq:= 19607843;
			when 154=> freq:= 19480519;
			when 155=> freq:= 19354838;
			when 156=> freq:= 19230769;
			when 157=> freq:= 19108280;
			when 158=> freq:= 18987341;
			when 159=> freq:= 18867924;
			when 160=> freq:= 18750000;
			when 161=> freq:= 18633540;
			when 162=> freq:= 18518518;
			when 163=> freq:= 18404908;
			when 164=> freq:= 18292682;
			when 165=> freq:= 18181818;
			when 166=> freq:= 18072289;
			when 167=> freq:= 17964071;
			when 168=> freq:= 17857142;
			when 169=> freq:= 17751479;
			when 170=> freq:= 17647058;
			when 171=> freq:= 17543859;
			when 172=> freq:= 17441860;
			when 173=> freq:= 17341040;
			when 174=> freq:= 17241379;
			when 175=> freq:= 17142857;
			when 176=> freq:= 17045454;
			when 177=> freq:= 16949152;
			when 178=> freq:= 16853932;
			when 179=> freq:= 16759776;
			when 180=> freq:= 16666666;
			when 181=> freq:= 16574585;
			when 182=> freq:= 16483516;
			when 183=> freq:= 16393442;
			when 184=> freq:= 16304347;
			when 185=> freq:= 16216216;
			when 186=> freq:= 16129032;
			when 187=> freq:= 16042780;
			when 188=> freq:= 15957446;
			when 189=> freq:= 15873015;
			when 190=> freq:= 15789473;
			when 191=> freq:= 15706806;
			when 192=> freq:= 15625000;
			when 193=> freq:= 15544041;
			when 194=> freq:= 15463917;
			when 195=> freq:= 15384615;
			when 196=> freq:= 15306122;
			when 197=> freq:= 15228426;
			when 198=> freq:= 15151515;
			when 199=> freq:= 15075376;
			when 200=> freq:= 15000000;
			when 201=> freq:= 14925373;
			when 202=> freq:= 14851485;
			when 203=> freq:= 14778325;
			when 204=> freq:= 14705882;
			when 205=> freq:= 14634146;
			when 206=> freq:= 14563106;
			when 207=> freq:= 14492753;
			when 208=> freq:= 14423076;
			when 209=> freq:= 14354067;
			when 210=> freq:= 14285714;
			when 211=> freq:= 14218009;
			when 212=> freq:= 14150943;
			when 213=> freq:= 14084507;
			when 214=> freq:= 14018691;
			when 215=> freq:= 13953488;
			when 216=> freq:= 13888888;
			when 217=> freq:= 13824884;
			when 218=> freq:= 13761467;
			when 219=> freq:= 13698630;
			when 220=> freq:= 13636363;
			when 221=> freq:= 13574660;
			when 222=> freq:= 13513513;
			when 223=> freq:= 13452914;
			when 224=> freq:= 13392857;
			when 225=> freq:= 13333333;
			when 226=> freq:= 13274336;
			when 227=> freq:= 13215859;
			when 228=> freq:= 13157894;
			when 229=> freq:= 13100436;
			when 230=> freq:= 13043478;
			when 231=> freq:= 12987013;
			when 232=> freq:= 12931034;
			when 233=> freq:= 12875536;
			when 234=> freq:= 12820512;
			when 235=> freq:= 12765957;
			when 236=> freq:= 12711864;
			when 237=> freq:= 12658227;
			when 238=> freq:= 12605042;
			when 239=> freq:= 12552301;
			when 240=> freq:= 12500000;
			when 241=> freq:= 12448132;
			when 242=> freq:= 12396694;
			when 243=> freq:= 12345679;
			when 244=> freq:= 12295082;
			when 245=> freq:= 12244898;
			when 246=> freq:= 12195122;
			when 247=> freq:= 12145749;
			when 248=> freq:= 12096774;
			when 249=> freq:= 12048192;
			when 250=> freq:= 12000000;
			when 251=> freq:= 11952191;
			when 252=> freq:= 11904761;
			when 253=> freq:= 11857707;
			when 254=> freq:= 11811023;
			when 255=> freq:= 11764705;
			when 256=> freq:= 11718750;
			when 257=> freq:= 11673151;
			when 258=> freq:= 11627907;
			when 259=> freq:= 11583011;
			when 260=> freq:= 11538461;
			when others => freq:= 50000000;
		end case;
	end if;
end process;

process(Clk, Resetn)
begin
	if Resetn='0' then counter<= (others=>'0');
	elsif (Clk' event and Clk = '0') then
		if counter < std_logic_vector(to_unsigned(freq -1,27)) then
			counter <= counter + 1;
		else
			counter <=(others=>'0');
		end if;
	end if;
end process;

process(counter)
begin
	if (counter >= freq/4-1 and counter < freq/2-1) then Secuencia_leds<="010";
	elsif (counter >= freq/2-1 and counter < freq*3/4-1) then Secuencia_leds<="011";
	elsif (counter >= freq*3/4-1 and counter < freq-1) then Secuencia_leds<="100";
	else Secuencia_leds<="001";
	end if;
end process;

process(Compas)
begin
	case Compas is
		when "0001" =>
			if (counter= freq-1 or counter< t_10ms -1) then Secuencia_sonido<= '1';
			else Secuencia_sonido<= '0';
			end if; 
		when "0010" => 
			if (counter= freq-1 or counter< t_10ms -1) then Secuencia_sonido<= '1';
			elsif (counter>= freq/2-1 and counter< freq/2 +t_10ms -1) then Secuencia_sonido<= '1';
			else Secuencia_sonido<= '0';
			end if;
		when "0011" =>
			if (counter= freq-1 or counter < t_10ms-1) then Secuencia_sonido<= '1';
			elsif (counter>=freq/3-1 and counter < freq/3 + t_10ms - 1) then Secuencia_sonido<= '1';
			elsif (counter>=freq*2/3-1 and counter < freq*2/3 + t_10ms -1) then Secuencia_sonido<= '1';
			else Secuencia_sonido<= '0';
			end if;
		when "0100" => 
			if (counter=freq-1 or counter< t_10ms-1) then Secuencia_sonido<= '1';
			elsif (counter>=freq/4-1 and counter<freq/4 + t_10ms -1) then Secuencia_sonido<= '1';
			elsif (counter>=freq/2-1 and counter<freq/2 + t_10ms -1) then Secuencia_sonido<= '1';
			elsif (counter>=freq*3/4-1  and counter<freq*3/4 + t_10ms -1) then Secuencia_sonido<= '1';
			else Secuencia_sonido<= '0';
			end if;
		when others =>
	end case;	
end process;
end Solucion;